`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/12/2022 12:47:17 PM
// Design Name: 
// Module Name: NbitSLT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NbitSLT #(parameter N = 32)(
    output [N-1:0] outval, 
    input [N-1:0] R2, 
    input [N-1:0] R3,
    input [N-1:0] inval //result of R2-R3
    );
    
    
    
endmodule
